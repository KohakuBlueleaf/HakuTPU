module DSP # (
    parameter integer INPUTREG = 1,
    parameter integer OUTPUTREG = 1,
    parameter integer DSPPIPEREG = 1,
    parameter integer CONTROLREG = 1,
    parameter integer NEEDPREADDER = 1
)(
    input clk,
    input rst,
    input enable,
    input signed [29:0] A,
    input signed [17:0] B,
    input signed [47:0] C,
    input signed [26:0] D,
    input signed [47:0] PCIN,
    input [8:0] OPMODE,
    input [4:0] INMODE,
    input [3:0] ALUMODE,
    output signed [47:0] P,
    output signed [47:0] PCOUT,
    output signed [29:0] ACOUT,
    output signed [17:0] BCOUT
);
    DSP48E2 #(
        .AMULTSEL(NEEDPREADDER ? "AD" : "A"),
        .AREG(INPUTREG),
        .ACASCREG(INPUTREG),
        .BREG(INPUTREG),
        .BCASCREG(INPUTREG),
        .MREG(DSPPIPEREG),
        .ADREG(DSPPIPEREG),
        .CREG(INPUTREG),
        .DREG(INPUTREG),
        .PREG(OUTPUTREG),
        .INMODEREG(CONTROLREG),
        .OPMODEREG(CONTROLREG),
        .ALUMODEREG(CONTROLREG)
    ) dsp_unit (
        .RSTA(rst),
        .RSTALLCARRYIN(rst),
        .RSTALUMODE(rst),
        .RSTB(rst),
        .RSTC(rst),
        .RSTCTRL(rst),
        .RSTD(rst),
        .RSTINMODE(rst),
        .RSTM(rst),
        .RSTP(rst),
        .CEA1(enable),
        .CEA2(enable),
        .CEAD(enable),
        .CEALUMODE(enable),
        .CEB1(enable),
        .CEB2(enable),
        .CEC(enable),
        .CECARRYIN(enable),
        .CECTRL(enable),
        .CED(enable),
        .CEINMODE(enable),
        .CEM(enable),
        .CEP(enable),
        .A(A),
        .B(B),
        .C(C),
        .D(D),
        .PCIN(PCIN),
        .CLK(clk),
        .ALUMODE(ALUMODE),
        .INMODE(INMODE),
        .OPMODE(OPMODE), // (A+D) * B + C + PCIN
        .P(P),
        .PCOUT(PCOUT),
        .ACOUT(ACOUT),
        .BCOUT(BCOUT)
    );
endmodule