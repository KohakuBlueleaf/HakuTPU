module FP12Inverse (
    input [11:0] a,
    output reg [15:0] b
);
    // input FP12 (E5M6) a;
    // output FP16 (E5M10) 1/a;
    // implement by LUT6_2 directly
    // a = 2^e * 1.m, 1/a = 2^-e * 1/(1.m), where 1/(1.m) is 6bit input 10bit output
    // real_e = e-15, -real_e = (-e + 30) - 15, final_e = -e + 30
    // if e!=0, mantissa = 1.m, 1/1.m = (0.5, 1], which means we need shift in exponent
    // therefore, if e!=0 and mantissa!=0, we need to minus 1 in exponent
    // NOTE: in this module we didn't handled 1/inf and 1/NaN, 
    //       they should be handled by ALU design directly
    wire sign = a[11];
    wire [4:0] exp = a[10:6];
    wire [5:0] mant = a[5:0];
    wire [10:0] mant_out;
    wire [10:0] subnorm_out;

    MultiBitLut #(
        .input_bits(6),
        .output_bits(11),
        .INIT({
            64'b0000000000000000000000000000000000000000000000000000000000000001,
            64'b0000000000000000000000000000000000000000001111111111111111111110,
            64'b0000000000000000000000000111111111111111110000000000001111111110,
            64'b0000000000000011111111111000000000111111110000000111110000011110,
            64'b0000000111111100000011111000001111000011110000111000110001100110,
            64'b0001111000111100011100111000110011001100110011011011010010101010,
            64'b0110011001001101101101001011010101010101010101101101100111000000,
            64'b1010101010010110110110011001110000000000000111001001010100110000,
            64'b0000000111001100100101010101101110000000011001010011101110101000,
            64'b0000111001010101001100000011001001000000101011111010010010000100,
            64'b0001001011000000100010000101011100110011000010001001010000000000
        })
    ) mlut (
        .in(mant),
        .out(mant_out)
    );

    MultiBitLut #(
        .input_bits(6),
        .output_bits(11),
        .INIT({
            // if the msb output bit is 1 it means NaN, fill all 1
            64'b0000000000000000000000000000000111111111111111111111111111111111,
            64'b0000000000000000000001111111111111111111111111111111111111111111,
            64'b0000000000001111111110000001111111111111111111111111111111111111,
            64'b0000000111110000011110001110011111111111111111111111111111111111,
            64'b0001111000110001100110010010101111111111111111111111111111111111,
            64'b0110011011010010101010110110000111111111111111111111111111111111,
            64'b1010101101100111111111101101100111111111111111111111111111111111,
            64'b0000011011010110000001100111010111111111111111111111111111111111,
            64'b0001101001111101000010110101000111111111111111111111111111111111,
            64'b0010111101000100100000110010001111111111111111111111111111111111,
            64'b0100100000001111010100000110000111111111111111111111111111111111
        })
    ) mlut_subnorm (
        .in(mant),
        .out(subnorm_out)
    );

    always @(*) begin
        if(exp==5'b00000) begin
            b = {sign, 4'b1111, subnorm_out};
        end else if(exp==5'b11101) begin
            b = {sign, 6'b1, mant_out[9:1]};
        end else if (exp==5'b11110) begin
            b = {sign, 7'b1, mant_out[9:2]};
        end else begin
            b = {sign, -exp + 5'd29 + mant_out[10], mant_out[9:0]};
        end
    end
endmodule